



module registers_ctrl 
#(
    parameter C_WIDTH = 32
)
(
    input iwClk,
    input iwRst,

)
{
};

endmodule
